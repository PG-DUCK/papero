-- soc_system.vhd

-- Generated using ACDS version 20.1 711

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system is
	port (
		button_pio_external_connection_export  : in    std_logic_vector(3 downto 0)  := (others => '0'); -- button_pio_external_connection.export
		clk_clk                                : in    std_logic                     := '0';             --                            clk.clk
		dipsw_pio_external_connection_export   : in    std_logic_vector(9 downto 0)  := (others => '0'); --  dipsw_pio_external_connection.export
		fast_fifo_fpga_to_hps_clk_clk          : in    std_logic                     := '0';             --      fast_fifo_fpga_to_hps_clk.clk
		fast_fifo_fpga_to_hps_in_writedata     : in    std_logic_vector(31 downto 0) := (others => '0'); --       fast_fifo_fpga_to_hps_in.writedata
		fast_fifo_fpga_to_hps_in_write         : in    std_logic                     := '0';             --                               .write
		fast_fifo_fpga_to_hps_in_waitrequest   : out   std_logic;                                        --                               .waitrequest
		fast_fifo_fpga_to_hps_in_csr_address   : in    std_logic_vector(2 downto 0)  := (others => '0'); --   fast_fifo_fpga_to_hps_in_csr.address
		fast_fifo_fpga_to_hps_in_csr_read      : in    std_logic                     := '0';             --                               .read
		fast_fifo_fpga_to_hps_in_csr_writedata : in    std_logic_vector(31 downto 0) := (others => '0'); --                               .writedata
		fast_fifo_fpga_to_hps_in_csr_write     : in    std_logic                     := '0';             --                               .write
		fast_fifo_fpga_to_hps_in_csr_readdata  : out   std_logic_vector(31 downto 0);                    --                               .readdata
		fast_fifo_fpga_to_hps_rst_reset_n      : in    std_logic                     := '0';             --      fast_fifo_fpga_to_hps_rst.reset_n
		fifo_fpga_to_hps_clk_clk               : in    std_logic                     := '0';             --           fifo_fpga_to_hps_clk.clk
		fifo_fpga_to_hps_in_writedata          : in    std_logic_vector(31 downto 0) := (others => '0'); --            fifo_fpga_to_hps_in.writedata
		fifo_fpga_to_hps_in_write              : in    std_logic                     := '0';             --                               .write
		fifo_fpga_to_hps_in_waitrequest        : out   std_logic;                                        --                               .waitrequest
		fifo_fpga_to_hps_in_csr_address        : in    std_logic_vector(2 downto 0)  := (others => '0'); --        fifo_fpga_to_hps_in_csr.address
		fifo_fpga_to_hps_in_csr_read           : in    std_logic                     := '0';             --                               .read
		fifo_fpga_to_hps_in_csr_writedata      : in    std_logic_vector(31 downto 0) := (others => '0'); --                               .writedata
		fifo_fpga_to_hps_in_csr_write          : in    std_logic                     := '0';             --                               .write
		fifo_fpga_to_hps_in_csr_readdata       : out   std_logic_vector(31 downto 0);                    --                               .readdata
		fifo_fpga_to_hps_rst_reset_n           : in    std_logic                     := '0';             --           fifo_fpga_to_hps_rst.reset_n
		fifo_hps_to_fpga_clk_clk               : in    std_logic                     := '0';             --           fifo_hps_to_fpga_clk.clk
		fifo_hps_to_fpga_out_readdata          : out   std_logic_vector(31 downto 0);                    --           fifo_hps_to_fpga_out.readdata
		fifo_hps_to_fpga_out_read              : in    std_logic                     := '0';             --                               .read
		fifo_hps_to_fpga_out_waitrequest       : out   std_logic;                                        --                               .waitrequest
		fifo_hps_to_fpga_out_csr_address       : in    std_logic_vector(2 downto 0)  := (others => '0'); --       fifo_hps_to_fpga_out_csr.address
		fifo_hps_to_fpga_out_csr_read          : in    std_logic                     := '0';             --                               .read
		fifo_hps_to_fpga_out_csr_writedata     : in    std_logic_vector(31 downto 0) := (others => '0'); --                               .writedata
		fifo_hps_to_fpga_out_csr_write         : in    std_logic                     := '0';             --                               .write
		fifo_hps_to_fpga_out_csr_readdata      : out   std_logic_vector(31 downto 0);                    --                               .readdata
		fifo_hps_to_fpga_rst_reset_n           : in    std_logic                     := '0';             --           fifo_hps_to_fpga_rst.reset_n
		hps_0_f2h_cold_reset_req_reset_n       : in    std_logic                     := '0';             --       hps_0_f2h_cold_reset_req.reset_n
		hps_0_f2h_debug_reset_req_reset_n      : in    std_logic                     := '0';             --      hps_0_f2h_debug_reset_req.reset_n
		hps_0_f2h_stm_hw_events_stm_hwevents   : in    std_logic_vector(27 downto 0) := (others => '0'); --        hps_0_f2h_stm_hw_events.stm_hwevents
		hps_0_f2h_warm_reset_req_reset_n       : in    std_logic                     := '0';             --       hps_0_f2h_warm_reset_req.reset_n
		hps_0_h2f_reset_reset_n                : out   std_logic;                                        --                hps_0_h2f_reset.reset_n
		hps_0_h2f_user0_clock_clk              : out   std_logic;                                        --          hps_0_h2f_user0_clock.clk
		hps_0_h2f_user1_clock_clk              : out   std_logic;                                        --          hps_0_h2f_user1_clock.clk
		hps_0_hps_io_hps_io_emac1_inst_TX_CLK  : out   std_logic;                                        --                   hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		hps_0_hps_io_hps_io_emac1_inst_TXD0    : out   std_logic;                                        --                               .hps_io_emac1_inst_TXD0
		hps_0_hps_io_hps_io_emac1_inst_TXD1    : out   std_logic;                                        --                               .hps_io_emac1_inst_TXD1
		hps_0_hps_io_hps_io_emac1_inst_TXD2    : out   std_logic;                                        --                               .hps_io_emac1_inst_TXD2
		hps_0_hps_io_hps_io_emac1_inst_TXD3    : out   std_logic;                                        --                               .hps_io_emac1_inst_TXD3
		hps_0_hps_io_hps_io_emac1_inst_RXD0    : in    std_logic                     := '0';             --                               .hps_io_emac1_inst_RXD0
		hps_0_hps_io_hps_io_emac1_inst_MDIO    : inout std_logic                     := '0';             --                               .hps_io_emac1_inst_MDIO
		hps_0_hps_io_hps_io_emac1_inst_MDC     : out   std_logic;                                        --                               .hps_io_emac1_inst_MDC
		hps_0_hps_io_hps_io_emac1_inst_RX_CTL  : in    std_logic                     := '0';             --                               .hps_io_emac1_inst_RX_CTL
		hps_0_hps_io_hps_io_emac1_inst_TX_CTL  : out   std_logic;                                        --                               .hps_io_emac1_inst_TX_CTL
		hps_0_hps_io_hps_io_emac1_inst_RX_CLK  : in    std_logic                     := '0';             --                               .hps_io_emac1_inst_RX_CLK
		hps_0_hps_io_hps_io_emac1_inst_RXD1    : in    std_logic                     := '0';             --                               .hps_io_emac1_inst_RXD1
		hps_0_hps_io_hps_io_emac1_inst_RXD2    : in    std_logic                     := '0';             --                               .hps_io_emac1_inst_RXD2
		hps_0_hps_io_hps_io_emac1_inst_RXD3    : in    std_logic                     := '0';             --                               .hps_io_emac1_inst_RXD3
		hps_0_hps_io_hps_io_qspi_inst_IO0      : inout std_logic                     := '0';             --                               .hps_io_qspi_inst_IO0
		hps_0_hps_io_hps_io_qspi_inst_IO1      : inout std_logic                     := '0';             --                               .hps_io_qspi_inst_IO1
		hps_0_hps_io_hps_io_qspi_inst_IO2      : inout std_logic                     := '0';             --                               .hps_io_qspi_inst_IO2
		hps_0_hps_io_hps_io_qspi_inst_IO3      : inout std_logic                     := '0';             --                               .hps_io_qspi_inst_IO3
		hps_0_hps_io_hps_io_qspi_inst_SS0      : out   std_logic;                                        --                               .hps_io_qspi_inst_SS0
		hps_0_hps_io_hps_io_qspi_inst_CLK      : out   std_logic;                                        --                               .hps_io_qspi_inst_CLK
		hps_0_hps_io_hps_io_sdio_inst_CMD      : inout std_logic                     := '0';             --                               .hps_io_sdio_inst_CMD
		hps_0_hps_io_hps_io_sdio_inst_D0       : inout std_logic                     := '0';             --                               .hps_io_sdio_inst_D0
		hps_0_hps_io_hps_io_sdio_inst_D1       : inout std_logic                     := '0';             --                               .hps_io_sdio_inst_D1
		hps_0_hps_io_hps_io_sdio_inst_CLK      : out   std_logic;                                        --                               .hps_io_sdio_inst_CLK
		hps_0_hps_io_hps_io_sdio_inst_D2       : inout std_logic                     := '0';             --                               .hps_io_sdio_inst_D2
		hps_0_hps_io_hps_io_sdio_inst_D3       : inout std_logic                     := '0';             --                               .hps_io_sdio_inst_D3
		hps_0_hps_io_hps_io_usb1_inst_D0       : inout std_logic                     := '0';             --                               .hps_io_usb1_inst_D0
		hps_0_hps_io_hps_io_usb1_inst_D1       : inout std_logic                     := '0';             --                               .hps_io_usb1_inst_D1
		hps_0_hps_io_hps_io_usb1_inst_D2       : inout std_logic                     := '0';             --                               .hps_io_usb1_inst_D2
		hps_0_hps_io_hps_io_usb1_inst_D3       : inout std_logic                     := '0';             --                               .hps_io_usb1_inst_D3
		hps_0_hps_io_hps_io_usb1_inst_D4       : inout std_logic                     := '0';             --                               .hps_io_usb1_inst_D4
		hps_0_hps_io_hps_io_usb1_inst_D5       : inout std_logic                     := '0';             --                               .hps_io_usb1_inst_D5
		hps_0_hps_io_hps_io_usb1_inst_D6       : inout std_logic                     := '0';             --                               .hps_io_usb1_inst_D6
		hps_0_hps_io_hps_io_usb1_inst_D7       : inout std_logic                     := '0';             --                               .hps_io_usb1_inst_D7
		hps_0_hps_io_hps_io_usb1_inst_CLK      : in    std_logic                     := '0';             --                               .hps_io_usb1_inst_CLK
		hps_0_hps_io_hps_io_usb1_inst_STP      : out   std_logic;                                        --                               .hps_io_usb1_inst_STP
		hps_0_hps_io_hps_io_usb1_inst_DIR      : in    std_logic                     := '0';             --                               .hps_io_usb1_inst_DIR
		hps_0_hps_io_hps_io_usb1_inst_NXT      : in    std_logic                     := '0';             --                               .hps_io_usb1_inst_NXT
		hps_0_hps_io_hps_io_spim0_inst_CLK     : out   std_logic;                                        --                               .hps_io_spim0_inst_CLK
		hps_0_hps_io_hps_io_spim0_inst_MOSI    : out   std_logic;                                        --                               .hps_io_spim0_inst_MOSI
		hps_0_hps_io_hps_io_spim0_inst_MISO    : in    std_logic                     := '0';             --                               .hps_io_spim0_inst_MISO
		hps_0_hps_io_hps_io_spim0_inst_SS0     : out   std_logic;                                        --                               .hps_io_spim0_inst_SS0
		hps_0_hps_io_hps_io_spim1_inst_CLK     : out   std_logic;                                        --                               .hps_io_spim1_inst_CLK
		hps_0_hps_io_hps_io_spim1_inst_MOSI    : out   std_logic;                                        --                               .hps_io_spim1_inst_MOSI
		hps_0_hps_io_hps_io_spim1_inst_MISO    : in    std_logic                     := '0';             --                               .hps_io_spim1_inst_MISO
		hps_0_hps_io_hps_io_spim1_inst_SS0     : out   std_logic;                                        --                               .hps_io_spim1_inst_SS0
		hps_0_hps_io_hps_io_uart0_inst_RX      : in    std_logic                     := '0';             --                               .hps_io_uart0_inst_RX
		hps_0_hps_io_hps_io_uart0_inst_TX      : out   std_logic;                                        --                               .hps_io_uart0_inst_TX
		hps_0_hps_io_hps_io_i2c0_inst_SDA      : inout std_logic                     := '0';             --                               .hps_io_i2c0_inst_SDA
		hps_0_hps_io_hps_io_i2c0_inst_SCL      : inout std_logic                     := '0';             --                               .hps_io_i2c0_inst_SCL
		hps_0_hps_io_hps_io_i2c1_inst_SDA      : inout std_logic                     := '0';             --                               .hps_io_i2c1_inst_SDA
		hps_0_hps_io_hps_io_i2c1_inst_SCL      : inout std_logic                     := '0';             --                               .hps_io_i2c1_inst_SCL
		hps_0_hps_io_hps_io_gpio_inst_GPIO09   : inout std_logic                     := '0';             --                               .hps_io_gpio_inst_GPIO09
		hps_0_hps_io_hps_io_gpio_inst_GPIO35   : inout std_logic                     := '0';             --                               .hps_io_gpio_inst_GPIO35
		hps_0_hps_io_hps_io_gpio_inst_GPIO37   : inout std_logic                     := '0';             --                               .hps_io_gpio_inst_GPIO37
		hps_0_hps_io_hps_io_gpio_inst_GPIO40   : inout std_logic                     := '0';             --                               .hps_io_gpio_inst_GPIO40
		hps_0_hps_io_hps_io_gpio_inst_GPIO41   : inout std_logic                     := '0';             --                               .hps_io_gpio_inst_GPIO41
		hps_0_hps_io_hps_io_gpio_inst_GPIO44   : inout std_logic                     := '0';             --                               .hps_io_gpio_inst_GPIO44
		hps_0_hps_io_hps_io_gpio_inst_GPIO48   : inout std_logic                     := '0';             --                               .hps_io_gpio_inst_GPIO48
		hps_0_hps_io_hps_io_gpio_inst_GPIO53   : inout std_logic                     := '0';             --                               .hps_io_gpio_inst_GPIO53
		hps_0_hps_io_hps_io_gpio_inst_GPIO54   : inout std_logic                     := '0';             --                               .hps_io_gpio_inst_GPIO54
		hps_0_hps_io_hps_io_gpio_inst_GPIO61   : inout std_logic                     := '0';             --                               .hps_io_gpio_inst_GPIO61
		led_pio_external_connection_export     : out   std_logic_vector(9 downto 0);                     --    led_pio_external_connection.export
		memory_mem_a                           : out   std_logic_vector(14 downto 0);                    --                         memory.mem_a
		memory_mem_ba                          : out   std_logic_vector(2 downto 0);                     --                               .mem_ba
		memory_mem_ck                          : out   std_logic;                                        --                               .mem_ck
		memory_mem_ck_n                        : out   std_logic;                                        --                               .mem_ck_n
		memory_mem_cke                         : out   std_logic;                                        --                               .mem_cke
		memory_mem_cs_n                        : out   std_logic;                                        --                               .mem_cs_n
		memory_mem_ras_n                       : out   std_logic;                                        --                               .mem_ras_n
		memory_mem_cas_n                       : out   std_logic;                                        --                               .mem_cas_n
		memory_mem_we_n                        : out   std_logic;                                        --                               .mem_we_n
		memory_mem_reset_n                     : out   std_logic;                                        --                               .mem_reset_n
		memory_mem_dq                          : inout std_logic_vector(31 downto 0) := (others => '0'); --                               .mem_dq
		memory_mem_dqs                         : inout std_logic_vector(3 downto 0)  := (others => '0'); --                               .mem_dqs
		memory_mem_dqs_n                       : inout std_logic_vector(3 downto 0)  := (others => '0'); --                               .mem_dqs_n
		memory_mem_odt                         : out   std_logic;                                        --                               .mem_odt
		memory_mem_dm                          : out   std_logic_vector(3 downto 0);                     --                               .mem_dm
		memory_oct_rzqin                       : in    std_logic                     := '0';             --                               .oct_rzqin
		regaddr_pio_export                     : out   std_logic_vector(31 downto 0);                    --                    regaddr_pio.export
		regcontent_pio_export                  : in    std_logic_vector(31 downto 0) := (others => '0'); --                 regcontent_pio.export
		reset_reset_n                          : in    std_logic                     := '0'              --                          reset.reset_n
	);
end entity soc_system;

architecture rtl of soc_system is
	component soc_system_RegAddr_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component soc_system_RegAddr_pio;

	component soc_system_RegContent_pio is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component soc_system_RegContent_pio;

	component soc_system_button_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component soc_system_button_pio;

	component soc_system_dipsw_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component soc_system_dipsw_pio;

	component soc_system_fast_fifo_FPGA_to_HPS is
		port (
			wrclock                          : in  std_logic                     := 'X';             -- clk
			wrreset_n                        : in  std_logic                     := 'X';             -- reset_n
			rdclock                          : in  std_logic                     := 'X';             -- clk
			rdreset_n                        : in  std_logic                     := 'X';             -- reset_n
			avalonmm_write_slave_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalonmm_write_slave_write       : in  std_logic                     := 'X';             -- write
			avalonmm_write_slave_waitrequest : out std_logic;                                        -- waitrequest
			avalonmm_read_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			avalonmm_read_slave_read         : in  std_logic                     := 'X';             -- read
			avalonmm_read_slave_waitrequest  : out std_logic;                                        -- waitrequest
			rdclk_control_slave_address      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			rdclk_control_slave_read         : in  std_logic                     := 'X';             -- read
			rdclk_control_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			rdclk_control_slave_write        : in  std_logic                     := 'X';             -- write
			rdclk_control_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			wrclk_control_slave_address      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			wrclk_control_slave_read         : in  std_logic                     := 'X';             -- read
			wrclk_control_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			wrclk_control_slave_write        : in  std_logic                     := 'X';             -- write
			wrclk_control_slave_readdata     : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component soc_system_fast_fifo_FPGA_to_HPS;

	component soc_system_fifo_FPGA_to_HPS is
		port (
			wrclock                          : in  std_logic                     := 'X';             -- clk
			wrreset_n                        : in  std_logic                     := 'X';             -- reset_n
			rdclock                          : in  std_logic                     := 'X';             -- clk
			rdreset_n                        : in  std_logic                     := 'X';             -- reset_n
			avalonmm_write_slave_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalonmm_write_slave_write       : in  std_logic                     := 'X';             -- write
			avalonmm_write_slave_waitrequest : out std_logic;                                        -- waitrequest
			avalonmm_read_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			avalonmm_read_slave_read         : in  std_logic                     := 'X';             -- read
			avalonmm_read_slave_waitrequest  : out std_logic;                                        -- waitrequest
			rdclk_control_slave_address      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			rdclk_control_slave_read         : in  std_logic                     := 'X';             -- read
			rdclk_control_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			rdclk_control_slave_write        : in  std_logic                     := 'X';             -- write
			rdclk_control_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			wrclk_control_slave_address      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			wrclk_control_slave_read         : in  std_logic                     := 'X';             -- read
			wrclk_control_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			wrclk_control_slave_write        : in  std_logic                     := 'X';             -- write
			wrclk_control_slave_readdata     : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component soc_system_fifo_FPGA_to_HPS;

	component soc_system_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			f2h_cold_rst_req_n       : in    std_logic                      := 'X';             -- reset_n
			f2h_dbg_rst_req_n        : in    std_logic                      := 'X';             -- reset_n
			f2h_warm_rst_req_n       : in    std_logic                      := 'X';             -- reset_n
			h2f_user0_clk            : out   std_logic;                                         -- clk
			h2f_user1_clk            : out   std_logic;                                         -- clk
			f2h_stm_hwevents         : in    std_logic_vector(27 downto 0)  := (others => 'X'); -- stm_hwevents
			mem_a                    : out   std_logic_vector(14 downto 0);                     -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                      -- mem_ba
			mem_ck                   : out   std_logic;                                         -- mem_ck
			mem_ck_n                 : out   std_logic;                                         -- mem_ck_n
			mem_cke                  : out   std_logic;                                         -- mem_cke
			mem_cs_n                 : out   std_logic;                                         -- mem_cs_n
			mem_ras_n                : out   std_logic;                                         -- mem_ras_n
			mem_cas_n                : out   std_logic;                                         -- mem_cas_n
			mem_we_n                 : out   std_logic;                                         -- mem_we_n
			mem_reset_n              : out   std_logic;                                         -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                         -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                      -- mem_dm
			oct_rzqin                : in    std_logic                      := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                         -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                         -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                         -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                         -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                         -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                      := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                         -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                         -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_qspi_inst_IO0     : inout std_logic                      := 'X';             -- hps_io_qspi_inst_IO0
			hps_io_qspi_inst_IO1     : inout std_logic                      := 'X';             -- hps_io_qspi_inst_IO1
			hps_io_qspi_inst_IO2     : inout std_logic                      := 'X';             -- hps_io_qspi_inst_IO2
			hps_io_qspi_inst_IO3     : inout std_logic                      := 'X';             -- hps_io_qspi_inst_IO3
			hps_io_qspi_inst_SS0     : out   std_logic;                                         -- hps_io_qspi_inst_SS0
			hps_io_qspi_inst_CLK     : out   std_logic;                                         -- hps_io_qspi_inst_CLK
			hps_io_sdio_inst_CMD     : inout std_logic                      := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                         -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     : out   std_logic;                                         -- hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_spim0_inst_CLK    : out   std_logic;                                         -- hps_io_spim0_inst_CLK
			hps_io_spim0_inst_MOSI   : out   std_logic;                                         -- hps_io_spim0_inst_MOSI
			hps_io_spim0_inst_MISO   : in    std_logic                      := 'X';             -- hps_io_spim0_inst_MISO
			hps_io_spim0_inst_SS0    : out   std_logic;                                         -- hps_io_spim0_inst_SS0
			hps_io_spim1_inst_CLK    : out   std_logic;                                         -- hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   : out   std_logic;                                         -- hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   : in    std_logic                      := 'X';             -- hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    : out   std_logic;                                         -- hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     : in    std_logic                      := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                         -- hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     : inout std_logic                      := 'X';             -- hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     : inout std_logic                      := 'X';             -- hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     : inout std_logic                      := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     : inout std_logic                      := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO37  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO37
			hps_io_gpio_inst_GPIO40  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO41  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO41
			hps_io_gpio_inst_GPIO44  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO44
			hps_io_gpio_inst_GPIO48  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO61
			h2f_rst_n                : out   std_logic;                                         -- reset_n
			f2h_sdram0_clk           : in    std_logic                      := 'X';             -- clk
			f2h_sdram0_ADDRESS       : in    std_logic_vector(26 downto 0)  := (others => 'X'); -- address
			f2h_sdram0_BURSTCOUNT    : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- burstcount
			f2h_sdram0_WAITREQUEST   : out   std_logic;                                         -- waitrequest
			f2h_sdram0_READDATA      : out   std_logic_vector(255 downto 0);                    -- readdata
			f2h_sdram0_READDATAVALID : out   std_logic;                                         -- readdatavalid
			f2h_sdram0_READ          : in    std_logic                      := 'X';             -- read
			f2h_sdram0_WRITEDATA     : in    std_logic_vector(255 downto 0) := (others => 'X'); -- writedata
			f2h_sdram0_BYTEENABLE    : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- byteenable
			f2h_sdram0_WRITE         : in    std_logic                      := 'X';             -- write
			h2f_axi_clk              : in    std_logic                      := 'X';             -- clk
			h2f_AWID                 : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_AWADDR               : out   std_logic_vector(29 downto 0);                     -- awaddr
			h2f_AWLEN                : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_AWSIZE               : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_AWBURST              : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_AWLOCK               : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_AWCACHE              : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_AWPROT               : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_AWVALID              : out   std_logic;                                         -- awvalid
			h2f_AWREADY              : in    std_logic                      := 'X';             -- awready
			h2f_WID                  : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_WDATA                : out   std_logic_vector(63 downto 0);                     -- wdata
			h2f_WSTRB                : out   std_logic_vector(7 downto 0);                      -- wstrb
			h2f_WLAST                : out   std_logic;                                         -- wlast
			h2f_WVALID               : out   std_logic;                                         -- wvalid
			h2f_WREADY               : in    std_logic                      := 'X';             -- wready
			h2f_BID                  : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_BRESP                : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_BVALID               : in    std_logic                      := 'X';             -- bvalid
			h2f_BREADY               : out   std_logic;                                         -- bready
			h2f_ARID                 : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_ARADDR               : out   std_logic_vector(29 downto 0);                     -- araddr
			h2f_ARLEN                : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_ARSIZE               : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_ARBURST              : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_ARLOCK               : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_ARCACHE              : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_ARPROT               : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_ARVALID              : out   std_logic;                                         -- arvalid
			h2f_ARREADY              : in    std_logic                      := 'X';             -- arready
			h2f_RID                  : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_RDATA                : in    std_logic_vector(63 downto 0)  := (others => 'X'); -- rdata
			h2f_RRESP                : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_RLAST                : in    std_logic                      := 'X';             -- rlast
			h2f_RVALID               : in    std_logic                      := 'X';             -- rvalid
			h2f_RREADY               : out   std_logic;                                         -- rready
			f2h_axi_clk              : in    std_logic                      := 'X';             -- clk
			f2h_AWID                 : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- awid
			f2h_AWADDR               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- awaddr
			f2h_AWLEN                : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			f2h_AWSIZE               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			f2h_AWBURST              : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			f2h_AWLOCK               : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			f2h_AWCACHE              : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			f2h_AWPROT               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			f2h_AWVALID              : in    std_logic                      := 'X';             -- awvalid
			f2h_AWREADY              : out   std_logic;                                         -- awready
			f2h_AWUSER               : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- awuser
			f2h_WID                  : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- wid
			f2h_WDATA                : in    std_logic_vector(63 downto 0)  := (others => 'X'); -- wdata
			f2h_WSTRB                : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- wstrb
			f2h_WLAST                : in    std_logic                      := 'X';             -- wlast
			f2h_WVALID               : in    std_logic                      := 'X';             -- wvalid
			f2h_WREADY               : out   std_logic;                                         -- wready
			f2h_BID                  : out   std_logic_vector(7 downto 0);                      -- bid
			f2h_BRESP                : out   std_logic_vector(1 downto 0);                      -- bresp
			f2h_BVALID               : out   std_logic;                                         -- bvalid
			f2h_BREADY               : in    std_logic                      := 'X';             -- bready
			f2h_ARID                 : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- arid
			f2h_ARADDR               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- araddr
			f2h_ARLEN                : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			f2h_ARSIZE               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			f2h_ARBURST              : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			f2h_ARLOCK               : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			f2h_ARCACHE              : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			f2h_ARPROT               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			f2h_ARVALID              : in    std_logic                      := 'X';             -- arvalid
			f2h_ARREADY              : out   std_logic;                                         -- arready
			f2h_ARUSER               : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- aruser
			f2h_RID                  : out   std_logic_vector(7 downto 0);                      -- rid
			f2h_RDATA                : out   std_logic_vector(63 downto 0);                     -- rdata
			f2h_RRESP                : out   std_logic_vector(1 downto 0);                      -- rresp
			f2h_RLAST                : out   std_logic;                                         -- rlast
			f2h_RVALID               : out   std_logic;                                         -- rvalid
			f2h_RREADY               : in    std_logic                      := 'X';             -- rready
			h2f_lw_axi_clk           : in    std_logic                      := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                     -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                         -- awvalid
			h2f_lw_AWREADY           : in    std_logic                      := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                     -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                      -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                         -- wlast
			h2f_lw_WVALID            : out   std_logic;                                         -- wvalid
			h2f_lw_WREADY            : in    std_logic                      := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                      := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                         -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                     -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                         -- arvalid
			h2f_lw_ARREADY           : in    std_logic                      := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                      := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                      := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic;                                         -- rready
			f2h_irq_p0               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- irq
			f2h_irq_p1               : in    std_logic_vector(31 downto 0)  := (others => 'X')  -- irq
		);
	end component soc_system_hps_0;

	component soc_system_led_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component soc_system_led_pio;

	component altera_avalon_mm_bridge is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			HDL_ADDR_WIDTH    : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(14 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic;                                        -- debugaccess
			s0_response      : out std_logic_vector(1 downto 0);                     -- response
			m0_response      : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- response
		);
	end component altera_avalon_mm_bridge;

	component soc_system_sysid_qsys is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component soc_system_sysid_qsys;

	component soc_system_mm_interconnect_0 is
		port (
			hps_0_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_0_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			hps_0_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_0_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_0_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_0_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_0_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_0_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_0_h2f_lw_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_0_h2f_lw_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_0_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_0_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_0_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_0_h2f_lw_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_0_h2f_lw_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_0_h2f_lw_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_0_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_0_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_0_h2f_lw_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_0_h2f_lw_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_0_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_0_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			hps_0_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_0_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_0_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_0_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_0_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_0_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_0_h2f_lw_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_0_h2f_lw_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_0_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_0_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                    -- rdata
			hps_0_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_0_h2f_lw_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_0_h2f_lw_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_0_h2f_lw_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			clk_0_clk_clk                                                       : in  std_logic                     := 'X';             -- clk
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			mm_bridge_0_reset_reset_bridge_in_reset_reset                       : in  std_logic                     := 'X';             -- reset
			mm_bridge_0_s0_address                                              : out std_logic_vector(14 downto 0);                    -- address
			mm_bridge_0_s0_write                                                : out std_logic;                                        -- write
			mm_bridge_0_s0_read                                                 : out std_logic;                                        -- read
			mm_bridge_0_s0_readdata                                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mm_bridge_0_s0_writedata                                            : out std_logic_vector(31 downto 0);                    -- writedata
			mm_bridge_0_s0_burstcount                                           : out std_logic_vector(0 downto 0);                     -- burstcount
			mm_bridge_0_s0_byteenable                                           : out std_logic_vector(3 downto 0);                     -- byteenable
			mm_bridge_0_s0_readdatavalid                                        : in  std_logic                     := 'X';             -- readdatavalid
			mm_bridge_0_s0_waitrequest                                          : in  std_logic                     := 'X';             -- waitrequest
			mm_bridge_0_s0_debugaccess                                          : out std_logic                                         -- debugaccess
		);
	end component soc_system_mm_interconnect_0;

	component soc_system_mm_interconnect_1 is
		port (
			clk_0_clk_clk                                 : in  std_logic                     := 'X';             -- clk
			mm_bridge_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			mm_bridge_0_m0_address                        : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			mm_bridge_0_m0_waitrequest                    : out std_logic;                                        -- waitrequest
			mm_bridge_0_m0_burstcount                     : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			mm_bridge_0_m0_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			mm_bridge_0_m0_read                           : in  std_logic                     := 'X';             -- read
			mm_bridge_0_m0_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			mm_bridge_0_m0_readdatavalid                  : out std_logic;                                        -- readdatavalid
			mm_bridge_0_m0_write                          : in  std_logic                     := 'X';             -- write
			mm_bridge_0_m0_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			mm_bridge_0_m0_debugaccess                    : in  std_logic                     := 'X';             -- debugaccess
			button_pio_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			button_pio_s1_write                           : out std_logic;                                        -- write
			button_pio_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			button_pio_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			button_pio_s1_chipselect                      : out std_logic;                                        -- chipselect
			dipsw_pio_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			dipsw_pio_s1_write                            : out std_logic;                                        -- write
			dipsw_pio_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			dipsw_pio_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			dipsw_pio_s1_chipselect                       : out std_logic;                                        -- chipselect
			fast_fifo_FPGA_to_HPS_out_read                : out std_logic;                                        -- read
			fast_fifo_FPGA_to_HPS_out_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fast_fifo_FPGA_to_HPS_out_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			fast_fifo_FPGA_to_HPS_out_csr_address         : out std_logic_vector(2 downto 0);                     -- address
			fast_fifo_FPGA_to_HPS_out_csr_write           : out std_logic;                                        -- write
			fast_fifo_FPGA_to_HPS_out_csr_read            : out std_logic;                                        -- read
			fast_fifo_FPGA_to_HPS_out_csr_readdata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fast_fifo_FPGA_to_HPS_out_csr_writedata       : out std_logic_vector(31 downto 0);                    -- writedata
			fifo_FPGA_to_HPS_out_read                     : out std_logic;                                        -- read
			fifo_FPGA_to_HPS_out_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fifo_FPGA_to_HPS_out_waitrequest              : in  std_logic                     := 'X';             -- waitrequest
			fifo_FPGA_to_HPS_out_csr_address              : out std_logic_vector(2 downto 0);                     -- address
			fifo_FPGA_to_HPS_out_csr_write                : out std_logic;                                        -- write
			fifo_FPGA_to_HPS_out_csr_read                 : out std_logic;                                        -- read
			fifo_FPGA_to_HPS_out_csr_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fifo_FPGA_to_HPS_out_csr_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			fifo_HPS_to_FPGA_in_write                     : out std_logic;                                        -- write
			fifo_HPS_to_FPGA_in_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			fifo_HPS_to_FPGA_in_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			fifo_HPS_to_FPGA_in_csr_address               : out std_logic_vector(2 downto 0);                     -- address
			fifo_HPS_to_FPGA_in_csr_write                 : out std_logic;                                        -- write
			fifo_HPS_to_FPGA_in_csr_read                  : out std_logic;                                        -- read
			fifo_HPS_to_FPGA_in_csr_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fifo_HPS_to_FPGA_in_csr_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			led_pio_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			led_pio_s1_write                              : out std_logic;                                        -- write
			led_pio_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_pio_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			led_pio_s1_chipselect                         : out std_logic;                                        -- chipselect
			RegAddr_pio_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			RegAddr_pio_s1_write                          : out std_logic;                                        -- write
			RegAddr_pio_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			RegAddr_pio_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			RegAddr_pio_s1_chipselect                     : out std_logic;                                        -- chipselect
			RegContent_pio_s1_address                     : out std_logic_vector(1 downto 0);                     -- address
			RegContent_pio_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sysid_qsys_control_slave_address              : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_control_slave_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component soc_system_mm_interconnect_1;

	component soc_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component soc_system_irq_mapper;

	component soc_system_irq_mapper_001 is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component soc_system_irq_mapper_001;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal hps_0_h2f_reset_reset                                     : std_logic;                     -- hps_0:h2f_rst_n -> [hps_0_h2f_reset_reset_n, hps_0_h2f_reset_reset_n:in]
	signal hps_0_h2f_lw_axi_master_awburst                           : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	signal hps_0_h2f_lw_axi_master_arlen                             : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	signal hps_0_h2f_lw_axi_master_wstrb                             : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	signal hps_0_h2f_lw_axi_master_wready                            : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	signal hps_0_h2f_lw_axi_master_rid                               : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	signal hps_0_h2f_lw_axi_master_rready                            : std_logic;                     -- hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	signal hps_0_h2f_lw_axi_master_awlen                             : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	signal hps_0_h2f_lw_axi_master_wid                               : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	signal hps_0_h2f_lw_axi_master_arcache                           : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	signal hps_0_h2f_lw_axi_master_wvalid                            : std_logic;                     -- hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	signal hps_0_h2f_lw_axi_master_araddr                            : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	signal hps_0_h2f_lw_axi_master_arprot                            : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	signal hps_0_h2f_lw_axi_master_awprot                            : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	signal hps_0_h2f_lw_axi_master_wdata                             : std_logic_vector(31 downto 0); -- hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	signal hps_0_h2f_lw_axi_master_arvalid                           : std_logic;                     -- hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	signal hps_0_h2f_lw_axi_master_awcache                           : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	signal hps_0_h2f_lw_axi_master_arid                              : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	signal hps_0_h2f_lw_axi_master_arlock                            : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	signal hps_0_h2f_lw_axi_master_awlock                            : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	signal hps_0_h2f_lw_axi_master_awaddr                            : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	signal hps_0_h2f_lw_axi_master_bresp                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	signal hps_0_h2f_lw_axi_master_arready                           : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	signal hps_0_h2f_lw_axi_master_rdata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	signal hps_0_h2f_lw_axi_master_awready                           : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	signal hps_0_h2f_lw_axi_master_arburst                           : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	signal hps_0_h2f_lw_axi_master_arsize                            : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	signal hps_0_h2f_lw_axi_master_bready                            : std_logic;                     -- hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	signal hps_0_h2f_lw_axi_master_rlast                             : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	signal hps_0_h2f_lw_axi_master_wlast                             : std_logic;                     -- hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	signal hps_0_h2f_lw_axi_master_rresp                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	signal hps_0_h2f_lw_axi_master_awid                              : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	signal hps_0_h2f_lw_axi_master_bid                               : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	signal hps_0_h2f_lw_axi_master_bvalid                            : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	signal hps_0_h2f_lw_axi_master_awsize                            : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	signal hps_0_h2f_lw_axi_master_awvalid                           : std_logic;                     -- hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	signal hps_0_h2f_lw_axi_master_rvalid                            : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	signal mm_interconnect_0_mm_bridge_0_s0_readdata                 : std_logic_vector(31 downto 0); -- mm_bridge_0:s0_readdata -> mm_interconnect_0:mm_bridge_0_s0_readdata
	signal mm_interconnect_0_mm_bridge_0_s0_waitrequest              : std_logic;                     -- mm_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_bridge_0_s0_waitrequest
	signal mm_interconnect_0_mm_bridge_0_s0_debugaccess              : std_logic;                     -- mm_interconnect_0:mm_bridge_0_s0_debugaccess -> mm_bridge_0:s0_debugaccess
	signal mm_interconnect_0_mm_bridge_0_s0_address                  : std_logic_vector(14 downto 0); -- mm_interconnect_0:mm_bridge_0_s0_address -> mm_bridge_0:s0_address
	signal mm_interconnect_0_mm_bridge_0_s0_read                     : std_logic;                     -- mm_interconnect_0:mm_bridge_0_s0_read -> mm_bridge_0:s0_read
	signal mm_interconnect_0_mm_bridge_0_s0_byteenable               : std_logic_vector(3 downto 0);  -- mm_interconnect_0:mm_bridge_0_s0_byteenable -> mm_bridge_0:s0_byteenable
	signal mm_interconnect_0_mm_bridge_0_s0_readdatavalid            : std_logic;                     -- mm_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_bridge_0_s0_readdatavalid
	signal mm_interconnect_0_mm_bridge_0_s0_write                    : std_logic;                     -- mm_interconnect_0:mm_bridge_0_s0_write -> mm_bridge_0:s0_write
	signal mm_interconnect_0_mm_bridge_0_s0_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:mm_bridge_0_s0_writedata -> mm_bridge_0:s0_writedata
	signal mm_interconnect_0_mm_bridge_0_s0_burstcount               : std_logic_vector(0 downto 0);  -- mm_interconnect_0:mm_bridge_0_s0_burstcount -> mm_bridge_0:s0_burstcount
	signal mm_bridge_0_m0_waitrequest                                : std_logic;                     -- mm_interconnect_1:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	signal mm_bridge_0_m0_readdata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_1:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	signal mm_bridge_0_m0_debugaccess                                : std_logic;                     -- mm_bridge_0:m0_debugaccess -> mm_interconnect_1:mm_bridge_0_m0_debugaccess
	signal mm_bridge_0_m0_address                                    : std_logic_vector(14 downto 0); -- mm_bridge_0:m0_address -> mm_interconnect_1:mm_bridge_0_m0_address
	signal mm_bridge_0_m0_read                                       : std_logic;                     -- mm_bridge_0:m0_read -> mm_interconnect_1:mm_bridge_0_m0_read
	signal mm_bridge_0_m0_byteenable                                 : std_logic_vector(3 downto 0);  -- mm_bridge_0:m0_byteenable -> mm_interconnect_1:mm_bridge_0_m0_byteenable
	signal mm_bridge_0_m0_readdatavalid                              : std_logic;                     -- mm_interconnect_1:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	signal mm_bridge_0_m0_writedata                                  : std_logic_vector(31 downto 0); -- mm_bridge_0:m0_writedata -> mm_interconnect_1:mm_bridge_0_m0_writedata
	signal mm_bridge_0_m0_write                                      : std_logic;                     -- mm_bridge_0:m0_write -> mm_interconnect_1:mm_bridge_0_m0_write
	signal mm_bridge_0_m0_burstcount                                 : std_logic_vector(0 downto 0);  -- mm_bridge_0:m0_burstcount -> mm_interconnect_1:mm_bridge_0_m0_burstcount
	signal mm_interconnect_1_sysid_qsys_control_slave_readdata       : std_logic_vector(31 downto 0); -- sysid_qsys:readdata -> mm_interconnect_1:sysid_qsys_control_slave_readdata
	signal mm_interconnect_1_sysid_qsys_control_slave_address        : std_logic_vector(0 downto 0);  -- mm_interconnect_1:sysid_qsys_control_slave_address -> sysid_qsys:address
	signal mm_interconnect_1_fifo_hps_to_fpga_in_waitrequest         : std_logic;                     -- fifo_HPS_to_FPGA:avalonmm_write_slave_waitrequest -> mm_interconnect_1:fifo_HPS_to_FPGA_in_waitrequest
	signal mm_interconnect_1_fifo_hps_to_fpga_in_write               : std_logic;                     -- mm_interconnect_1:fifo_HPS_to_FPGA_in_write -> fifo_HPS_to_FPGA:avalonmm_write_slave_write
	signal mm_interconnect_1_fifo_hps_to_fpga_in_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_1:fifo_HPS_to_FPGA_in_writedata -> fifo_HPS_to_FPGA:avalonmm_write_slave_writedata
	signal mm_interconnect_1_fifo_hps_to_fpga_in_csr_readdata        : std_logic_vector(31 downto 0); -- fifo_HPS_to_FPGA:wrclk_control_slave_readdata -> mm_interconnect_1:fifo_HPS_to_FPGA_in_csr_readdata
	signal mm_interconnect_1_fifo_hps_to_fpga_in_csr_address         : std_logic_vector(2 downto 0);  -- mm_interconnect_1:fifo_HPS_to_FPGA_in_csr_address -> fifo_HPS_to_FPGA:wrclk_control_slave_address
	signal mm_interconnect_1_fifo_hps_to_fpga_in_csr_read            : std_logic;                     -- mm_interconnect_1:fifo_HPS_to_FPGA_in_csr_read -> fifo_HPS_to_FPGA:wrclk_control_slave_read
	signal mm_interconnect_1_fifo_hps_to_fpga_in_csr_write           : std_logic;                     -- mm_interconnect_1:fifo_HPS_to_FPGA_in_csr_write -> fifo_HPS_to_FPGA:wrclk_control_slave_write
	signal mm_interconnect_1_fifo_hps_to_fpga_in_csr_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_1:fifo_HPS_to_FPGA_in_csr_writedata -> fifo_HPS_to_FPGA:wrclk_control_slave_writedata
	signal mm_interconnect_1_fifo_fpga_to_hps_out_readdata           : std_logic_vector(31 downto 0); -- fifo_FPGA_to_HPS:avalonmm_read_slave_readdata -> mm_interconnect_1:fifo_FPGA_to_HPS_out_readdata
	signal mm_interconnect_1_fifo_fpga_to_hps_out_waitrequest        : std_logic;                     -- fifo_FPGA_to_HPS:avalonmm_read_slave_waitrequest -> mm_interconnect_1:fifo_FPGA_to_HPS_out_waitrequest
	signal mm_interconnect_1_fifo_fpga_to_hps_out_read               : std_logic;                     -- mm_interconnect_1:fifo_FPGA_to_HPS_out_read -> fifo_FPGA_to_HPS:avalonmm_read_slave_read
	signal mm_interconnect_1_fast_fifo_fpga_to_hps_out_readdata      : std_logic_vector(31 downto 0); -- fast_fifo_FPGA_to_HPS:avalonmm_read_slave_readdata -> mm_interconnect_1:fast_fifo_FPGA_to_HPS_out_readdata
	signal mm_interconnect_1_fast_fifo_fpga_to_hps_out_waitrequest   : std_logic;                     -- fast_fifo_FPGA_to_HPS:avalonmm_read_slave_waitrequest -> mm_interconnect_1:fast_fifo_FPGA_to_HPS_out_waitrequest
	signal mm_interconnect_1_fast_fifo_fpga_to_hps_out_read          : std_logic;                     -- mm_interconnect_1:fast_fifo_FPGA_to_HPS_out_read -> fast_fifo_FPGA_to_HPS:avalonmm_read_slave_read
	signal mm_interconnect_1_fifo_fpga_to_hps_out_csr_readdata       : std_logic_vector(31 downto 0); -- fifo_FPGA_to_HPS:rdclk_control_slave_readdata -> mm_interconnect_1:fifo_FPGA_to_HPS_out_csr_readdata
	signal mm_interconnect_1_fifo_fpga_to_hps_out_csr_address        : std_logic_vector(2 downto 0);  -- mm_interconnect_1:fifo_FPGA_to_HPS_out_csr_address -> fifo_FPGA_to_HPS:rdclk_control_slave_address
	signal mm_interconnect_1_fifo_fpga_to_hps_out_csr_read           : std_logic;                     -- mm_interconnect_1:fifo_FPGA_to_HPS_out_csr_read -> fifo_FPGA_to_HPS:rdclk_control_slave_read
	signal mm_interconnect_1_fifo_fpga_to_hps_out_csr_write          : std_logic;                     -- mm_interconnect_1:fifo_FPGA_to_HPS_out_csr_write -> fifo_FPGA_to_HPS:rdclk_control_slave_write
	signal mm_interconnect_1_fifo_fpga_to_hps_out_csr_writedata      : std_logic_vector(31 downto 0); -- mm_interconnect_1:fifo_FPGA_to_HPS_out_csr_writedata -> fifo_FPGA_to_HPS:rdclk_control_slave_writedata
	signal mm_interconnect_1_fast_fifo_fpga_to_hps_out_csr_readdata  : std_logic_vector(31 downto 0); -- fast_fifo_FPGA_to_HPS:rdclk_control_slave_readdata -> mm_interconnect_1:fast_fifo_FPGA_to_HPS_out_csr_readdata
	signal mm_interconnect_1_fast_fifo_fpga_to_hps_out_csr_address   : std_logic_vector(2 downto 0);  -- mm_interconnect_1:fast_fifo_FPGA_to_HPS_out_csr_address -> fast_fifo_FPGA_to_HPS:rdclk_control_slave_address
	signal mm_interconnect_1_fast_fifo_fpga_to_hps_out_csr_read      : std_logic;                     -- mm_interconnect_1:fast_fifo_FPGA_to_HPS_out_csr_read -> fast_fifo_FPGA_to_HPS:rdclk_control_slave_read
	signal mm_interconnect_1_fast_fifo_fpga_to_hps_out_csr_write     : std_logic;                     -- mm_interconnect_1:fast_fifo_FPGA_to_HPS_out_csr_write -> fast_fifo_FPGA_to_HPS:rdclk_control_slave_write
	signal mm_interconnect_1_fast_fifo_fpga_to_hps_out_csr_writedata : std_logic_vector(31 downto 0); -- mm_interconnect_1:fast_fifo_FPGA_to_HPS_out_csr_writedata -> fast_fifo_FPGA_to_HPS:rdclk_control_slave_writedata
	signal mm_interconnect_1_button_pio_s1_chipselect                : std_logic;                     -- mm_interconnect_1:button_pio_s1_chipselect -> button_pio:chipselect
	signal mm_interconnect_1_button_pio_s1_readdata                  : std_logic_vector(31 downto 0); -- button_pio:readdata -> mm_interconnect_1:button_pio_s1_readdata
	signal mm_interconnect_1_button_pio_s1_address                   : std_logic_vector(1 downto 0);  -- mm_interconnect_1:button_pio_s1_address -> button_pio:address
	signal mm_interconnect_1_button_pio_s1_write                     : std_logic;                     -- mm_interconnect_1:button_pio_s1_write -> mm_interconnect_1_button_pio_s1_write:in
	signal mm_interconnect_1_button_pio_s1_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_1:button_pio_s1_writedata -> button_pio:writedata
	signal mm_interconnect_1_dipsw_pio_s1_chipselect                 : std_logic;                     -- mm_interconnect_1:dipsw_pio_s1_chipselect -> dipsw_pio:chipselect
	signal mm_interconnect_1_dipsw_pio_s1_readdata                   : std_logic_vector(31 downto 0); -- dipsw_pio:readdata -> mm_interconnect_1:dipsw_pio_s1_readdata
	signal mm_interconnect_1_dipsw_pio_s1_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_1:dipsw_pio_s1_address -> dipsw_pio:address
	signal mm_interconnect_1_dipsw_pio_s1_write                      : std_logic;                     -- mm_interconnect_1:dipsw_pio_s1_write -> mm_interconnect_1_dipsw_pio_s1_write:in
	signal mm_interconnect_1_dipsw_pio_s1_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_1:dipsw_pio_s1_writedata -> dipsw_pio:writedata
	signal mm_interconnect_1_led_pio_s1_chipselect                   : std_logic;                     -- mm_interconnect_1:led_pio_s1_chipselect -> led_pio:chipselect
	signal mm_interconnect_1_led_pio_s1_readdata                     : std_logic_vector(31 downto 0); -- led_pio:readdata -> mm_interconnect_1:led_pio_s1_readdata
	signal mm_interconnect_1_led_pio_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_1:led_pio_s1_address -> led_pio:address
	signal mm_interconnect_1_led_pio_s1_write                        : std_logic;                     -- mm_interconnect_1:led_pio_s1_write -> mm_interconnect_1_led_pio_s1_write:in
	signal mm_interconnect_1_led_pio_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_1:led_pio_s1_writedata -> led_pio:writedata
	signal mm_interconnect_1_regcontent_pio_s1_readdata              : std_logic_vector(31 downto 0); -- RegContent_pio:readdata -> mm_interconnect_1:RegContent_pio_s1_readdata
	signal mm_interconnect_1_regcontent_pio_s1_address               : std_logic_vector(1 downto 0);  -- mm_interconnect_1:RegContent_pio_s1_address -> RegContent_pio:address
	signal mm_interconnect_1_regaddr_pio_s1_chipselect               : std_logic;                     -- mm_interconnect_1:RegAddr_pio_s1_chipselect -> RegAddr_pio:chipselect
	signal mm_interconnect_1_regaddr_pio_s1_readdata                 : std_logic_vector(31 downto 0); -- RegAddr_pio:readdata -> mm_interconnect_1:RegAddr_pio_s1_readdata
	signal mm_interconnect_1_regaddr_pio_s1_address                  : std_logic_vector(1 downto 0);  -- mm_interconnect_1:RegAddr_pio_s1_address -> RegAddr_pio:address
	signal mm_interconnect_1_regaddr_pio_s1_write                    : std_logic;                     -- mm_interconnect_1:RegAddr_pio_s1_write -> mm_interconnect_1_regaddr_pio_s1_write:in
	signal mm_interconnect_1_regaddr_pio_s1_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_1:RegAddr_pio_s1_writedata -> RegAddr_pio:writedata
	signal irq_mapper_receiver0_irq                                  : std_logic;                     -- button_pio:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                  : std_logic;                     -- dipsw_pio:irq -> irq_mapper:receiver1_irq
	signal hps_0_f2h_irq0_irq                                        : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	signal hps_0_f2h_irq1_irq                                        : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	signal rst_controller_reset_out_reset                            : std_logic;                     -- rst_controller:reset_out -> [mm_bridge_0:reset, mm_interconnect_0:mm_bridge_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mm_bridge_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                        : std_logic;                     -- rst_controller_001:reset_out -> mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	signal hps_0_h2f_reset_reset_n_ports_inv                         : std_logic;                     -- hps_0_h2f_reset_reset_n:inv -> rst_controller_001:reset_in0
	signal reset_reset_n_ports_inv                                   : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_1_button_pio_s1_write_ports_inv           : std_logic;                     -- mm_interconnect_1_button_pio_s1_write:inv -> button_pio:write_n
	signal mm_interconnect_1_dipsw_pio_s1_write_ports_inv            : std_logic;                     -- mm_interconnect_1_dipsw_pio_s1_write:inv -> dipsw_pio:write_n
	signal mm_interconnect_1_led_pio_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_1_led_pio_s1_write:inv -> led_pio:write_n
	signal mm_interconnect_1_regaddr_pio_s1_write_ports_inv          : std_logic;                     -- mm_interconnect_1_regaddr_pio_s1_write:inv -> RegAddr_pio:write_n
	signal rst_controller_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_reset_out_reset:inv -> [RegAddr_pio:reset_n, RegContent_pio:reset_n, button_pio:reset_n, dipsw_pio:reset_n, fast_fifo_FPGA_to_HPS:rdreset_n, fifo_FPGA_to_HPS:rdreset_n, fifo_HPS_to_FPGA:wrreset_n, led_pio:reset_n, sysid_qsys:reset_n]

begin

	regaddr_pio : component soc_system_RegAddr_pio
		port map (
			clk        => clk_clk,                                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_1_regaddr_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_regaddr_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_regaddr_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_regaddr_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_regaddr_pio_s1_readdata,        --                    .readdata
			out_port   => regaddr_pio_export                                -- external_connection.export
		);

	regcontent_pio : component soc_system_RegContent_pio
		port map (
			clk      => clk_clk,                                      --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address  => mm_interconnect_1_regcontent_pio_s1_address,  --                  s1.address
			readdata => mm_interconnect_1_regcontent_pio_s1_readdata, --                    .readdata
			in_port  => regcontent_pio_export                         -- external_connection.export
		);

	button_pio : component soc_system_button_pio
		port map (
			clk        => clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_1_button_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_button_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_button_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_button_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_button_pio_s1_readdata,        --                    .readdata
			in_port    => button_pio_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver0_irq                         --                 irq.irq
		);

	dipsw_pio : component soc_system_dipsw_pio
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_1_dipsw_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_dipsw_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_dipsw_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_dipsw_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_dipsw_pio_s1_readdata,        --                    .readdata
			in_port    => dipsw_pio_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver1_irq                        --                 irq.irq
		);

	fast_fifo_fpga_to_hps : component soc_system_fast_fifo_FPGA_to_HPS
		port map (
			wrclock                          => fast_fifo_fpga_to_hps_clk_clk,                             --    clk_in.clk
			wrreset_n                        => fast_fifo_fpga_to_hps_rst_reset_n,                         --  reset_in.reset_n
			rdclock                          => clk_clk,                                                   --   clk_out.clk
			rdreset_n                        => rst_controller_reset_out_reset_ports_inv,                  -- reset_out.reset_n
			avalonmm_write_slave_writedata   => fast_fifo_fpga_to_hps_in_writedata,                        --        in.writedata
			avalonmm_write_slave_write       => fast_fifo_fpga_to_hps_in_write,                            --          .write
			avalonmm_write_slave_waitrequest => fast_fifo_fpga_to_hps_in_waitrequest,                      --          .waitrequest
			avalonmm_read_slave_readdata     => mm_interconnect_1_fast_fifo_fpga_to_hps_out_readdata,      --       out.readdata
			avalonmm_read_slave_read         => mm_interconnect_1_fast_fifo_fpga_to_hps_out_read,          --          .read
			avalonmm_read_slave_waitrequest  => mm_interconnect_1_fast_fifo_fpga_to_hps_out_waitrequest,   --          .waitrequest
			rdclk_control_slave_address      => mm_interconnect_1_fast_fifo_fpga_to_hps_out_csr_address,   --   out_csr.address
			rdclk_control_slave_read         => mm_interconnect_1_fast_fifo_fpga_to_hps_out_csr_read,      --          .read
			rdclk_control_slave_writedata    => mm_interconnect_1_fast_fifo_fpga_to_hps_out_csr_writedata, --          .writedata
			rdclk_control_slave_write        => mm_interconnect_1_fast_fifo_fpga_to_hps_out_csr_write,     --          .write
			rdclk_control_slave_readdata     => mm_interconnect_1_fast_fifo_fpga_to_hps_out_csr_readdata,  --          .readdata
			wrclk_control_slave_address      => fast_fifo_fpga_to_hps_in_csr_address,                      --    in_csr.address
			wrclk_control_slave_read         => fast_fifo_fpga_to_hps_in_csr_read,                         --          .read
			wrclk_control_slave_writedata    => fast_fifo_fpga_to_hps_in_csr_writedata,                    --          .writedata
			wrclk_control_slave_write        => fast_fifo_fpga_to_hps_in_csr_write,                        --          .write
			wrclk_control_slave_readdata     => fast_fifo_fpga_to_hps_in_csr_readdata                      --          .readdata
		);

	fifo_fpga_to_hps : component soc_system_fifo_FPGA_to_HPS
		port map (
			wrclock                          => fifo_fpga_to_hps_clk_clk,                             --    clk_in.clk
			wrreset_n                        => fifo_fpga_to_hps_rst_reset_n,                         --  reset_in.reset_n
			rdclock                          => clk_clk,                                              --   clk_out.clk
			rdreset_n                        => rst_controller_reset_out_reset_ports_inv,             -- reset_out.reset_n
			avalonmm_write_slave_writedata   => fifo_fpga_to_hps_in_writedata,                        --        in.writedata
			avalonmm_write_slave_write       => fifo_fpga_to_hps_in_write,                            --          .write
			avalonmm_write_slave_waitrequest => fifo_fpga_to_hps_in_waitrequest,                      --          .waitrequest
			avalonmm_read_slave_readdata     => mm_interconnect_1_fifo_fpga_to_hps_out_readdata,      --       out.readdata
			avalonmm_read_slave_read         => mm_interconnect_1_fifo_fpga_to_hps_out_read,          --          .read
			avalonmm_read_slave_waitrequest  => mm_interconnect_1_fifo_fpga_to_hps_out_waitrequest,   --          .waitrequest
			rdclk_control_slave_address      => mm_interconnect_1_fifo_fpga_to_hps_out_csr_address,   --   out_csr.address
			rdclk_control_slave_read         => mm_interconnect_1_fifo_fpga_to_hps_out_csr_read,      --          .read
			rdclk_control_slave_writedata    => mm_interconnect_1_fifo_fpga_to_hps_out_csr_writedata, --          .writedata
			rdclk_control_slave_write        => mm_interconnect_1_fifo_fpga_to_hps_out_csr_write,     --          .write
			rdclk_control_slave_readdata     => mm_interconnect_1_fifo_fpga_to_hps_out_csr_readdata,  --          .readdata
			wrclk_control_slave_address      => fifo_fpga_to_hps_in_csr_address,                      --    in_csr.address
			wrclk_control_slave_read         => fifo_fpga_to_hps_in_csr_read,                         --          .read
			wrclk_control_slave_writedata    => fifo_fpga_to_hps_in_csr_writedata,                    --          .writedata
			wrclk_control_slave_write        => fifo_fpga_to_hps_in_csr_write,                        --          .write
			wrclk_control_slave_readdata     => fifo_fpga_to_hps_in_csr_readdata                      --          .readdata
		);

	fifo_hps_to_fpga : component soc_system_fifo_FPGA_to_HPS
		port map (
			wrclock                          => clk_clk,                                             --    clk_in.clk
			wrreset_n                        => rst_controller_reset_out_reset_ports_inv,            --  reset_in.reset_n
			rdclock                          => fifo_hps_to_fpga_clk_clk,                            --   clk_out.clk
			rdreset_n                        => fifo_hps_to_fpga_rst_reset_n,                        -- reset_out.reset_n
			avalonmm_write_slave_writedata   => mm_interconnect_1_fifo_hps_to_fpga_in_writedata,     --        in.writedata
			avalonmm_write_slave_write       => mm_interconnect_1_fifo_hps_to_fpga_in_write,         --          .write
			avalonmm_write_slave_waitrequest => mm_interconnect_1_fifo_hps_to_fpga_in_waitrequest,   --          .waitrequest
			avalonmm_read_slave_readdata     => fifo_hps_to_fpga_out_readdata,                       --       out.readdata
			avalonmm_read_slave_read         => fifo_hps_to_fpga_out_read,                           --          .read
			avalonmm_read_slave_waitrequest  => fifo_hps_to_fpga_out_waitrequest,                    --          .waitrequest
			rdclk_control_slave_address      => fifo_hps_to_fpga_out_csr_address,                    --   out_csr.address
			rdclk_control_slave_read         => fifo_hps_to_fpga_out_csr_read,                       --          .read
			rdclk_control_slave_writedata    => fifo_hps_to_fpga_out_csr_writedata,                  --          .writedata
			rdclk_control_slave_write        => fifo_hps_to_fpga_out_csr_write,                      --          .write
			rdclk_control_slave_readdata     => fifo_hps_to_fpga_out_csr_readdata,                   --          .readdata
			wrclk_control_slave_address      => mm_interconnect_1_fifo_hps_to_fpga_in_csr_address,   --    in_csr.address
			wrclk_control_slave_read         => mm_interconnect_1_fifo_hps_to_fpga_in_csr_read,      --          .read
			wrclk_control_slave_writedata    => mm_interconnect_1_fifo_hps_to_fpga_in_csr_writedata, --          .writedata
			wrclk_control_slave_write        => mm_interconnect_1_fifo_hps_to_fpga_in_csr_write,     --          .write
			wrclk_control_slave_readdata     => mm_interconnect_1_fifo_hps_to_fpga_in_csr_readdata   --          .readdata
		);

	hps_0 : component soc_system_hps_0
		generic map (
			F2S_Width => 2,
			S2F_Width => 2
		)
		port map (
			f2h_cold_rst_req_n       => hps_0_f2h_cold_reset_req_reset_n,      --  f2h_cold_reset_req.reset_n
			f2h_dbg_rst_req_n        => hps_0_f2h_debug_reset_req_reset_n,     -- f2h_debug_reset_req.reset_n
			f2h_warm_rst_req_n       => hps_0_f2h_warm_reset_req_reset_n,      --  f2h_warm_reset_req.reset_n
			h2f_user0_clk            => hps_0_h2f_user0_clock_clk,             --     h2f_user0_clock.clk
			h2f_user1_clk            => hps_0_h2f_user1_clock_clk,             --     h2f_user1_clock.clk
			f2h_stm_hwevents         => hps_0_f2h_stm_hw_events_stm_hwevents,  --   f2h_stm_hw_events.stm_hwevents
			mem_a                    => memory_mem_a,                          --              memory.mem_a
			mem_ba                   => memory_mem_ba,                         --                    .mem_ba
			mem_ck                   => memory_mem_ck,                         --                    .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                       --                    .mem_ck_n
			mem_cke                  => memory_mem_cke,                        --                    .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                       --                    .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                      --                    .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                      --                    .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                       --                    .mem_we_n
			mem_reset_n              => memory_mem_reset_n,                    --                    .mem_reset_n
			mem_dq                   => memory_mem_dq,                         --                    .mem_dq
			mem_dqs                  => memory_mem_dqs,                        --                    .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                      --                    .mem_dqs_n
			mem_odt                  => memory_mem_odt,                        --                    .mem_odt
			mem_dm                   => memory_mem_dm,                         --                    .mem_dm
			oct_rzqin                => memory_oct_rzqin,                      --                    .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_0_hps_io_hps_io_emac1_inst_TX_CLK, --              hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_0_hps_io_hps_io_emac1_inst_TXD0,   --                    .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_0_hps_io_hps_io_emac1_inst_TXD1,   --                    .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_0_hps_io_hps_io_emac1_inst_TXD2,   --                    .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_0_hps_io_hps_io_emac1_inst_TXD3,   --                    .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_0_hps_io_hps_io_emac1_inst_RXD0,   --                    .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_0_hps_io_hps_io_emac1_inst_MDIO,   --                    .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_0_hps_io_hps_io_emac1_inst_MDC,    --                    .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_0_hps_io_hps_io_emac1_inst_RX_CTL, --                    .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_0_hps_io_hps_io_emac1_inst_TX_CTL, --                    .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_0_hps_io_hps_io_emac1_inst_RX_CLK, --                    .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_0_hps_io_hps_io_emac1_inst_RXD1,   --                    .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_0_hps_io_hps_io_emac1_inst_RXD2,   --                    .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_0_hps_io_hps_io_emac1_inst_RXD3,   --                    .hps_io_emac1_inst_RXD3
			hps_io_qspi_inst_IO0     => hps_0_hps_io_hps_io_qspi_inst_IO0,     --                    .hps_io_qspi_inst_IO0
			hps_io_qspi_inst_IO1     => hps_0_hps_io_hps_io_qspi_inst_IO1,     --                    .hps_io_qspi_inst_IO1
			hps_io_qspi_inst_IO2     => hps_0_hps_io_hps_io_qspi_inst_IO2,     --                    .hps_io_qspi_inst_IO2
			hps_io_qspi_inst_IO3     => hps_0_hps_io_hps_io_qspi_inst_IO3,     --                    .hps_io_qspi_inst_IO3
			hps_io_qspi_inst_SS0     => hps_0_hps_io_hps_io_qspi_inst_SS0,     --                    .hps_io_qspi_inst_SS0
			hps_io_qspi_inst_CLK     => hps_0_hps_io_hps_io_qspi_inst_CLK,     --                    .hps_io_qspi_inst_CLK
			hps_io_sdio_inst_CMD     => hps_0_hps_io_hps_io_sdio_inst_CMD,     --                    .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_0_hps_io_hps_io_sdio_inst_D0,      --                    .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_0_hps_io_hps_io_sdio_inst_D1,      --                    .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_0_hps_io_hps_io_sdio_inst_CLK,     --                    .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_0_hps_io_hps_io_sdio_inst_D2,      --                    .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_0_hps_io_hps_io_sdio_inst_D3,      --                    .hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      => hps_0_hps_io_hps_io_usb1_inst_D0,      --                    .hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      => hps_0_hps_io_hps_io_usb1_inst_D1,      --                    .hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      => hps_0_hps_io_hps_io_usb1_inst_D2,      --                    .hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      => hps_0_hps_io_hps_io_usb1_inst_D3,      --                    .hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      => hps_0_hps_io_hps_io_usb1_inst_D4,      --                    .hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      => hps_0_hps_io_hps_io_usb1_inst_D5,      --                    .hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      => hps_0_hps_io_hps_io_usb1_inst_D6,      --                    .hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      => hps_0_hps_io_hps_io_usb1_inst_D7,      --                    .hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     => hps_0_hps_io_hps_io_usb1_inst_CLK,     --                    .hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     => hps_0_hps_io_hps_io_usb1_inst_STP,     --                    .hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     => hps_0_hps_io_hps_io_usb1_inst_DIR,     --                    .hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     => hps_0_hps_io_hps_io_usb1_inst_NXT,     --                    .hps_io_usb1_inst_NXT
			hps_io_spim0_inst_CLK    => hps_0_hps_io_hps_io_spim0_inst_CLK,    --                    .hps_io_spim0_inst_CLK
			hps_io_spim0_inst_MOSI   => hps_0_hps_io_hps_io_spim0_inst_MOSI,   --                    .hps_io_spim0_inst_MOSI
			hps_io_spim0_inst_MISO   => hps_0_hps_io_hps_io_spim0_inst_MISO,   --                    .hps_io_spim0_inst_MISO
			hps_io_spim0_inst_SS0    => hps_0_hps_io_hps_io_spim0_inst_SS0,    --                    .hps_io_spim0_inst_SS0
			hps_io_spim1_inst_CLK    => hps_0_hps_io_hps_io_spim1_inst_CLK,    --                    .hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   => hps_0_hps_io_hps_io_spim1_inst_MOSI,   --                    .hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   => hps_0_hps_io_hps_io_spim1_inst_MISO,   --                    .hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    => hps_0_hps_io_hps_io_spim1_inst_SS0,    --                    .hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     => hps_0_hps_io_hps_io_uart0_inst_RX,     --                    .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_0_hps_io_hps_io_uart0_inst_TX,     --                    .hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     => hps_0_hps_io_hps_io_i2c0_inst_SDA,     --                    .hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     => hps_0_hps_io_hps_io_i2c0_inst_SCL,     --                    .hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     => hps_0_hps_io_hps_io_i2c1_inst_SDA,     --                    .hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     => hps_0_hps_io_hps_io_i2c1_inst_SCL,     --                    .hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  => hps_0_hps_io_hps_io_gpio_inst_GPIO09,  --                    .hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  => hps_0_hps_io_hps_io_gpio_inst_GPIO35,  --                    .hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO37  => hps_0_hps_io_hps_io_gpio_inst_GPIO37,  --                    .hps_io_gpio_inst_GPIO37
			hps_io_gpio_inst_GPIO40  => hps_0_hps_io_hps_io_gpio_inst_GPIO40,  --                    .hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO41  => hps_0_hps_io_hps_io_gpio_inst_GPIO41,  --                    .hps_io_gpio_inst_GPIO41
			hps_io_gpio_inst_GPIO44  => hps_0_hps_io_hps_io_gpio_inst_GPIO44,  --                    .hps_io_gpio_inst_GPIO44
			hps_io_gpio_inst_GPIO48  => hps_0_hps_io_hps_io_gpio_inst_GPIO48,  --                    .hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53  => hps_0_hps_io_hps_io_gpio_inst_GPIO53,  --                    .hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  => hps_0_hps_io_hps_io_gpio_inst_GPIO54,  --                    .hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  => hps_0_hps_io_hps_io_gpio_inst_GPIO61,  --                    .hps_io_gpio_inst_GPIO61
			h2f_rst_n                => hps_0_h2f_reset_reset,                 --           h2f_reset.reset_n
			f2h_sdram0_clk           => clk_clk,                               --    f2h_sdram0_clock.clk
			f2h_sdram0_ADDRESS       => open,                                  --     f2h_sdram0_data.address
			f2h_sdram0_BURSTCOUNT    => open,                                  --                    .burstcount
			f2h_sdram0_WAITREQUEST   => open,                                  --                    .waitrequest
			f2h_sdram0_READDATA      => open,                                  --                    .readdata
			f2h_sdram0_READDATAVALID => open,                                  --                    .readdatavalid
			f2h_sdram0_READ          => open,                                  --                    .read
			f2h_sdram0_WRITEDATA     => open,                                  --                    .writedata
			f2h_sdram0_BYTEENABLE    => open,                                  --                    .byteenable
			f2h_sdram0_WRITE         => open,                                  --                    .write
			h2f_axi_clk              => clk_clk,                               --       h2f_axi_clock.clk
			h2f_AWID                 => open,                                  --      h2f_axi_master.awid
			h2f_AWADDR               => open,                                  --                    .awaddr
			h2f_AWLEN                => open,                                  --                    .awlen
			h2f_AWSIZE               => open,                                  --                    .awsize
			h2f_AWBURST              => open,                                  --                    .awburst
			h2f_AWLOCK               => open,                                  --                    .awlock
			h2f_AWCACHE              => open,                                  --                    .awcache
			h2f_AWPROT               => open,                                  --                    .awprot
			h2f_AWVALID              => open,                                  --                    .awvalid
			h2f_AWREADY              => open,                                  --                    .awready
			h2f_WID                  => open,                                  --                    .wid
			h2f_WDATA                => open,                                  --                    .wdata
			h2f_WSTRB                => open,                                  --                    .wstrb
			h2f_WLAST                => open,                                  --                    .wlast
			h2f_WVALID               => open,                                  --                    .wvalid
			h2f_WREADY               => open,                                  --                    .wready
			h2f_BID                  => open,                                  --                    .bid
			h2f_BRESP                => open,                                  --                    .bresp
			h2f_BVALID               => open,                                  --                    .bvalid
			h2f_BREADY               => open,                                  --                    .bready
			h2f_ARID                 => open,                                  --                    .arid
			h2f_ARADDR               => open,                                  --                    .araddr
			h2f_ARLEN                => open,                                  --                    .arlen
			h2f_ARSIZE               => open,                                  --                    .arsize
			h2f_ARBURST              => open,                                  --                    .arburst
			h2f_ARLOCK               => open,                                  --                    .arlock
			h2f_ARCACHE              => open,                                  --                    .arcache
			h2f_ARPROT               => open,                                  --                    .arprot
			h2f_ARVALID              => open,                                  --                    .arvalid
			h2f_ARREADY              => open,                                  --                    .arready
			h2f_RID                  => open,                                  --                    .rid
			h2f_RDATA                => open,                                  --                    .rdata
			h2f_RRESP                => open,                                  --                    .rresp
			h2f_RLAST                => open,                                  --                    .rlast
			h2f_RVALID               => open,                                  --                    .rvalid
			h2f_RREADY               => open,                                  --                    .rready
			f2h_axi_clk              => clk_clk,                               --       f2h_axi_clock.clk
			f2h_AWID                 => open,                                  --       f2h_axi_slave.awid
			f2h_AWADDR               => open,                                  --                    .awaddr
			f2h_AWLEN                => open,                                  --                    .awlen
			f2h_AWSIZE               => open,                                  --                    .awsize
			f2h_AWBURST              => open,                                  --                    .awburst
			f2h_AWLOCK               => open,                                  --                    .awlock
			f2h_AWCACHE              => open,                                  --                    .awcache
			f2h_AWPROT               => open,                                  --                    .awprot
			f2h_AWVALID              => open,                                  --                    .awvalid
			f2h_AWREADY              => open,                                  --                    .awready
			f2h_AWUSER               => open,                                  --                    .awuser
			f2h_WID                  => open,                                  --                    .wid
			f2h_WDATA                => open,                                  --                    .wdata
			f2h_WSTRB                => open,                                  --                    .wstrb
			f2h_WLAST                => open,                                  --                    .wlast
			f2h_WVALID               => open,                                  --                    .wvalid
			f2h_WREADY               => open,                                  --                    .wready
			f2h_BID                  => open,                                  --                    .bid
			f2h_BRESP                => open,                                  --                    .bresp
			f2h_BVALID               => open,                                  --                    .bvalid
			f2h_BREADY               => open,                                  --                    .bready
			f2h_ARID                 => open,                                  --                    .arid
			f2h_ARADDR               => open,                                  --                    .araddr
			f2h_ARLEN                => open,                                  --                    .arlen
			f2h_ARSIZE               => open,                                  --                    .arsize
			f2h_ARBURST              => open,                                  --                    .arburst
			f2h_ARLOCK               => open,                                  --                    .arlock
			f2h_ARCACHE              => open,                                  --                    .arcache
			f2h_ARPROT               => open,                                  --                    .arprot
			f2h_ARVALID              => open,                                  --                    .arvalid
			f2h_ARREADY              => open,                                  --                    .arready
			f2h_ARUSER               => open,                                  --                    .aruser
			f2h_RID                  => open,                                  --                    .rid
			f2h_RDATA                => open,                                  --                    .rdata
			f2h_RRESP                => open,                                  --                    .rresp
			f2h_RLAST                => open,                                  --                    .rlast
			f2h_RVALID               => open,                                  --                    .rvalid
			f2h_RREADY               => open,                                  --                    .rready
			h2f_lw_axi_clk           => clk_clk,                               --    h2f_lw_axi_clock.clk
			h2f_lw_AWID              => hps_0_h2f_lw_axi_master_awid,          --   h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => hps_0_h2f_lw_axi_master_awaddr,        --                    .awaddr
			h2f_lw_AWLEN             => hps_0_h2f_lw_axi_master_awlen,         --                    .awlen
			h2f_lw_AWSIZE            => hps_0_h2f_lw_axi_master_awsize,        --                    .awsize
			h2f_lw_AWBURST           => hps_0_h2f_lw_axi_master_awburst,       --                    .awburst
			h2f_lw_AWLOCK            => hps_0_h2f_lw_axi_master_awlock,        --                    .awlock
			h2f_lw_AWCACHE           => hps_0_h2f_lw_axi_master_awcache,       --                    .awcache
			h2f_lw_AWPROT            => hps_0_h2f_lw_axi_master_awprot,        --                    .awprot
			h2f_lw_AWVALID           => hps_0_h2f_lw_axi_master_awvalid,       --                    .awvalid
			h2f_lw_AWREADY           => hps_0_h2f_lw_axi_master_awready,       --                    .awready
			h2f_lw_WID               => hps_0_h2f_lw_axi_master_wid,           --                    .wid
			h2f_lw_WDATA             => hps_0_h2f_lw_axi_master_wdata,         --                    .wdata
			h2f_lw_WSTRB             => hps_0_h2f_lw_axi_master_wstrb,         --                    .wstrb
			h2f_lw_WLAST             => hps_0_h2f_lw_axi_master_wlast,         --                    .wlast
			h2f_lw_WVALID            => hps_0_h2f_lw_axi_master_wvalid,        --                    .wvalid
			h2f_lw_WREADY            => hps_0_h2f_lw_axi_master_wready,        --                    .wready
			h2f_lw_BID               => hps_0_h2f_lw_axi_master_bid,           --                    .bid
			h2f_lw_BRESP             => hps_0_h2f_lw_axi_master_bresp,         --                    .bresp
			h2f_lw_BVALID            => hps_0_h2f_lw_axi_master_bvalid,        --                    .bvalid
			h2f_lw_BREADY            => hps_0_h2f_lw_axi_master_bready,        --                    .bready
			h2f_lw_ARID              => hps_0_h2f_lw_axi_master_arid,          --                    .arid
			h2f_lw_ARADDR            => hps_0_h2f_lw_axi_master_araddr,        --                    .araddr
			h2f_lw_ARLEN             => hps_0_h2f_lw_axi_master_arlen,         --                    .arlen
			h2f_lw_ARSIZE            => hps_0_h2f_lw_axi_master_arsize,        --                    .arsize
			h2f_lw_ARBURST           => hps_0_h2f_lw_axi_master_arburst,       --                    .arburst
			h2f_lw_ARLOCK            => hps_0_h2f_lw_axi_master_arlock,        --                    .arlock
			h2f_lw_ARCACHE           => hps_0_h2f_lw_axi_master_arcache,       --                    .arcache
			h2f_lw_ARPROT            => hps_0_h2f_lw_axi_master_arprot,        --                    .arprot
			h2f_lw_ARVALID           => hps_0_h2f_lw_axi_master_arvalid,       --                    .arvalid
			h2f_lw_ARREADY           => hps_0_h2f_lw_axi_master_arready,       --                    .arready
			h2f_lw_RID               => hps_0_h2f_lw_axi_master_rid,           --                    .rid
			h2f_lw_RDATA             => hps_0_h2f_lw_axi_master_rdata,         --                    .rdata
			h2f_lw_RRESP             => hps_0_h2f_lw_axi_master_rresp,         --                    .rresp
			h2f_lw_RLAST             => hps_0_h2f_lw_axi_master_rlast,         --                    .rlast
			h2f_lw_RVALID            => hps_0_h2f_lw_axi_master_rvalid,        --                    .rvalid
			h2f_lw_RREADY            => hps_0_h2f_lw_axi_master_rready,        --                    .rready
			f2h_irq_p0               => hps_0_f2h_irq0_irq,                    --            f2h_irq0.irq
			f2h_irq_p1               => hps_0_f2h_irq1_irq                     --            f2h_irq1.irq
		);

	led_pio : component soc_system_led_pio
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_1_led_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_led_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_led_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_led_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_led_pio_s1_readdata,        --                    .readdata
			out_port   => led_pio_external_connection_export            -- external_connection.export
		);

	mm_bridge_0 : component altera_avalon_mm_bridge
		generic map (
			DATA_WIDTH        => 32,
			SYMBOL_WIDTH      => 8,
			HDL_ADDR_WIDTH    => 15,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 1,
			PIPELINE_RESPONSE => 1
		)
		port map (
			clk              => clk_clk,                                        --   clk.clk
			reset            => rst_controller_reset_out_reset,                 -- reset.reset
			s0_waitrequest   => mm_interconnect_0_mm_bridge_0_s0_waitrequest,   --    s0.waitrequest
			s0_readdata      => mm_interconnect_0_mm_bridge_0_s0_readdata,      --      .readdata
			s0_readdatavalid => mm_interconnect_0_mm_bridge_0_s0_readdatavalid, --      .readdatavalid
			s0_burstcount    => mm_interconnect_0_mm_bridge_0_s0_burstcount,    --      .burstcount
			s0_writedata     => mm_interconnect_0_mm_bridge_0_s0_writedata,     --      .writedata
			s0_address       => mm_interconnect_0_mm_bridge_0_s0_address,       --      .address
			s0_write         => mm_interconnect_0_mm_bridge_0_s0_write,         --      .write
			s0_read          => mm_interconnect_0_mm_bridge_0_s0_read,          --      .read
			s0_byteenable    => mm_interconnect_0_mm_bridge_0_s0_byteenable,    --      .byteenable
			s0_debugaccess   => mm_interconnect_0_mm_bridge_0_s0_debugaccess,   --      .debugaccess
			m0_waitrequest   => mm_bridge_0_m0_waitrequest,                     --    m0.waitrequest
			m0_readdata      => mm_bridge_0_m0_readdata,                        --      .readdata
			m0_readdatavalid => mm_bridge_0_m0_readdatavalid,                   --      .readdatavalid
			m0_burstcount    => mm_bridge_0_m0_burstcount,                      --      .burstcount
			m0_writedata     => mm_bridge_0_m0_writedata,                       --      .writedata
			m0_address       => mm_bridge_0_m0_address,                         --      .address
			m0_write         => mm_bridge_0_m0_write,                           --      .write
			m0_read          => mm_bridge_0_m0_read,                            --      .read
			m0_byteenable    => mm_bridge_0_m0_byteenable,                      --      .byteenable
			m0_debugaccess   => mm_bridge_0_m0_debugaccess,                     --      .debugaccess
			s0_response      => open,                                           -- (terminated)
			m0_response      => "00"                                            -- (terminated)
		);

	sysid_qsys : component soc_system_sysid_qsys
		port map (
			clock    => clk_clk,                                               --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,              --         reset.reset_n
			readdata => mm_interconnect_1_sysid_qsys_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_1_sysid_qsys_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component soc_system_mm_interconnect_0
		port map (
			hps_0_h2f_lw_axi_master_awid                                        => hps_0_h2f_lw_axi_master_awid,                   --                                       hps_0_h2f_lw_axi_master.awid
			hps_0_h2f_lw_axi_master_awaddr                                      => hps_0_h2f_lw_axi_master_awaddr,                 --                                                              .awaddr
			hps_0_h2f_lw_axi_master_awlen                                       => hps_0_h2f_lw_axi_master_awlen,                  --                                                              .awlen
			hps_0_h2f_lw_axi_master_awsize                                      => hps_0_h2f_lw_axi_master_awsize,                 --                                                              .awsize
			hps_0_h2f_lw_axi_master_awburst                                     => hps_0_h2f_lw_axi_master_awburst,                --                                                              .awburst
			hps_0_h2f_lw_axi_master_awlock                                      => hps_0_h2f_lw_axi_master_awlock,                 --                                                              .awlock
			hps_0_h2f_lw_axi_master_awcache                                     => hps_0_h2f_lw_axi_master_awcache,                --                                                              .awcache
			hps_0_h2f_lw_axi_master_awprot                                      => hps_0_h2f_lw_axi_master_awprot,                 --                                                              .awprot
			hps_0_h2f_lw_axi_master_awvalid                                     => hps_0_h2f_lw_axi_master_awvalid,                --                                                              .awvalid
			hps_0_h2f_lw_axi_master_awready                                     => hps_0_h2f_lw_axi_master_awready,                --                                                              .awready
			hps_0_h2f_lw_axi_master_wid                                         => hps_0_h2f_lw_axi_master_wid,                    --                                                              .wid
			hps_0_h2f_lw_axi_master_wdata                                       => hps_0_h2f_lw_axi_master_wdata,                  --                                                              .wdata
			hps_0_h2f_lw_axi_master_wstrb                                       => hps_0_h2f_lw_axi_master_wstrb,                  --                                                              .wstrb
			hps_0_h2f_lw_axi_master_wlast                                       => hps_0_h2f_lw_axi_master_wlast,                  --                                                              .wlast
			hps_0_h2f_lw_axi_master_wvalid                                      => hps_0_h2f_lw_axi_master_wvalid,                 --                                                              .wvalid
			hps_0_h2f_lw_axi_master_wready                                      => hps_0_h2f_lw_axi_master_wready,                 --                                                              .wready
			hps_0_h2f_lw_axi_master_bid                                         => hps_0_h2f_lw_axi_master_bid,                    --                                                              .bid
			hps_0_h2f_lw_axi_master_bresp                                       => hps_0_h2f_lw_axi_master_bresp,                  --                                                              .bresp
			hps_0_h2f_lw_axi_master_bvalid                                      => hps_0_h2f_lw_axi_master_bvalid,                 --                                                              .bvalid
			hps_0_h2f_lw_axi_master_bready                                      => hps_0_h2f_lw_axi_master_bready,                 --                                                              .bready
			hps_0_h2f_lw_axi_master_arid                                        => hps_0_h2f_lw_axi_master_arid,                   --                                                              .arid
			hps_0_h2f_lw_axi_master_araddr                                      => hps_0_h2f_lw_axi_master_araddr,                 --                                                              .araddr
			hps_0_h2f_lw_axi_master_arlen                                       => hps_0_h2f_lw_axi_master_arlen,                  --                                                              .arlen
			hps_0_h2f_lw_axi_master_arsize                                      => hps_0_h2f_lw_axi_master_arsize,                 --                                                              .arsize
			hps_0_h2f_lw_axi_master_arburst                                     => hps_0_h2f_lw_axi_master_arburst,                --                                                              .arburst
			hps_0_h2f_lw_axi_master_arlock                                      => hps_0_h2f_lw_axi_master_arlock,                 --                                                              .arlock
			hps_0_h2f_lw_axi_master_arcache                                     => hps_0_h2f_lw_axi_master_arcache,                --                                                              .arcache
			hps_0_h2f_lw_axi_master_arprot                                      => hps_0_h2f_lw_axi_master_arprot,                 --                                                              .arprot
			hps_0_h2f_lw_axi_master_arvalid                                     => hps_0_h2f_lw_axi_master_arvalid,                --                                                              .arvalid
			hps_0_h2f_lw_axi_master_arready                                     => hps_0_h2f_lw_axi_master_arready,                --                                                              .arready
			hps_0_h2f_lw_axi_master_rid                                         => hps_0_h2f_lw_axi_master_rid,                    --                                                              .rid
			hps_0_h2f_lw_axi_master_rdata                                       => hps_0_h2f_lw_axi_master_rdata,                  --                                                              .rdata
			hps_0_h2f_lw_axi_master_rresp                                       => hps_0_h2f_lw_axi_master_rresp,                  --                                                              .rresp
			hps_0_h2f_lw_axi_master_rlast                                       => hps_0_h2f_lw_axi_master_rlast,                  --                                                              .rlast
			hps_0_h2f_lw_axi_master_rvalid                                      => hps_0_h2f_lw_axi_master_rvalid,                 --                                                              .rvalid
			hps_0_h2f_lw_axi_master_rready                                      => hps_0_h2f_lw_axi_master_rready,                 --                                                              .rready
			clk_0_clk_clk                                                       => clk_clk,                                        --                                                     clk_0_clk.clk
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,             -- hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			mm_bridge_0_reset_reset_bridge_in_reset_reset                       => rst_controller_reset_out_reset,                 --                       mm_bridge_0_reset_reset_bridge_in_reset.reset
			mm_bridge_0_s0_address                                              => mm_interconnect_0_mm_bridge_0_s0_address,       --                                                mm_bridge_0_s0.address
			mm_bridge_0_s0_write                                                => mm_interconnect_0_mm_bridge_0_s0_write,         --                                                              .write
			mm_bridge_0_s0_read                                                 => mm_interconnect_0_mm_bridge_0_s0_read,          --                                                              .read
			mm_bridge_0_s0_readdata                                             => mm_interconnect_0_mm_bridge_0_s0_readdata,      --                                                              .readdata
			mm_bridge_0_s0_writedata                                            => mm_interconnect_0_mm_bridge_0_s0_writedata,     --                                                              .writedata
			mm_bridge_0_s0_burstcount                                           => mm_interconnect_0_mm_bridge_0_s0_burstcount,    --                                                              .burstcount
			mm_bridge_0_s0_byteenable                                           => mm_interconnect_0_mm_bridge_0_s0_byteenable,    --                                                              .byteenable
			mm_bridge_0_s0_readdatavalid                                        => mm_interconnect_0_mm_bridge_0_s0_readdatavalid, --                                                              .readdatavalid
			mm_bridge_0_s0_waitrequest                                          => mm_interconnect_0_mm_bridge_0_s0_waitrequest,   --                                                              .waitrequest
			mm_bridge_0_s0_debugaccess                                          => mm_interconnect_0_mm_bridge_0_s0_debugaccess    --                                                              .debugaccess
		);

	mm_interconnect_1 : component soc_system_mm_interconnect_1
		port map (
			clk_0_clk_clk                                 => clk_clk,                                                   --                               clk_0_clk.clk
			mm_bridge_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                            -- mm_bridge_0_reset_reset_bridge_in_reset.reset
			mm_bridge_0_m0_address                        => mm_bridge_0_m0_address,                                    --                          mm_bridge_0_m0.address
			mm_bridge_0_m0_waitrequest                    => mm_bridge_0_m0_waitrequest,                                --                                        .waitrequest
			mm_bridge_0_m0_burstcount                     => mm_bridge_0_m0_burstcount,                                 --                                        .burstcount
			mm_bridge_0_m0_byteenable                     => mm_bridge_0_m0_byteenable,                                 --                                        .byteenable
			mm_bridge_0_m0_read                           => mm_bridge_0_m0_read,                                       --                                        .read
			mm_bridge_0_m0_readdata                       => mm_bridge_0_m0_readdata,                                   --                                        .readdata
			mm_bridge_0_m0_readdatavalid                  => mm_bridge_0_m0_readdatavalid,                              --                                        .readdatavalid
			mm_bridge_0_m0_write                          => mm_bridge_0_m0_write,                                      --                                        .write
			mm_bridge_0_m0_writedata                      => mm_bridge_0_m0_writedata,                                  --                                        .writedata
			mm_bridge_0_m0_debugaccess                    => mm_bridge_0_m0_debugaccess,                                --                                        .debugaccess
			button_pio_s1_address                         => mm_interconnect_1_button_pio_s1_address,                   --                           button_pio_s1.address
			button_pio_s1_write                           => mm_interconnect_1_button_pio_s1_write,                     --                                        .write
			button_pio_s1_readdata                        => mm_interconnect_1_button_pio_s1_readdata,                  --                                        .readdata
			button_pio_s1_writedata                       => mm_interconnect_1_button_pio_s1_writedata,                 --                                        .writedata
			button_pio_s1_chipselect                      => mm_interconnect_1_button_pio_s1_chipselect,                --                                        .chipselect
			dipsw_pio_s1_address                          => mm_interconnect_1_dipsw_pio_s1_address,                    --                            dipsw_pio_s1.address
			dipsw_pio_s1_write                            => mm_interconnect_1_dipsw_pio_s1_write,                      --                                        .write
			dipsw_pio_s1_readdata                         => mm_interconnect_1_dipsw_pio_s1_readdata,                   --                                        .readdata
			dipsw_pio_s1_writedata                        => mm_interconnect_1_dipsw_pio_s1_writedata,                  --                                        .writedata
			dipsw_pio_s1_chipselect                       => mm_interconnect_1_dipsw_pio_s1_chipselect,                 --                                        .chipselect
			fast_fifo_FPGA_to_HPS_out_read                => mm_interconnect_1_fast_fifo_fpga_to_hps_out_read,          --               fast_fifo_FPGA_to_HPS_out.read
			fast_fifo_FPGA_to_HPS_out_readdata            => mm_interconnect_1_fast_fifo_fpga_to_hps_out_readdata,      --                                        .readdata
			fast_fifo_FPGA_to_HPS_out_waitrequest         => mm_interconnect_1_fast_fifo_fpga_to_hps_out_waitrequest,   --                                        .waitrequest
			fast_fifo_FPGA_to_HPS_out_csr_address         => mm_interconnect_1_fast_fifo_fpga_to_hps_out_csr_address,   --           fast_fifo_FPGA_to_HPS_out_csr.address
			fast_fifo_FPGA_to_HPS_out_csr_write           => mm_interconnect_1_fast_fifo_fpga_to_hps_out_csr_write,     --                                        .write
			fast_fifo_FPGA_to_HPS_out_csr_read            => mm_interconnect_1_fast_fifo_fpga_to_hps_out_csr_read,      --                                        .read
			fast_fifo_FPGA_to_HPS_out_csr_readdata        => mm_interconnect_1_fast_fifo_fpga_to_hps_out_csr_readdata,  --                                        .readdata
			fast_fifo_FPGA_to_HPS_out_csr_writedata       => mm_interconnect_1_fast_fifo_fpga_to_hps_out_csr_writedata, --                                        .writedata
			fifo_FPGA_to_HPS_out_read                     => mm_interconnect_1_fifo_fpga_to_hps_out_read,               --                    fifo_FPGA_to_HPS_out.read
			fifo_FPGA_to_HPS_out_readdata                 => mm_interconnect_1_fifo_fpga_to_hps_out_readdata,           --                                        .readdata
			fifo_FPGA_to_HPS_out_waitrequest              => mm_interconnect_1_fifo_fpga_to_hps_out_waitrequest,        --                                        .waitrequest
			fifo_FPGA_to_HPS_out_csr_address              => mm_interconnect_1_fifo_fpga_to_hps_out_csr_address,        --                fifo_FPGA_to_HPS_out_csr.address
			fifo_FPGA_to_HPS_out_csr_write                => mm_interconnect_1_fifo_fpga_to_hps_out_csr_write,          --                                        .write
			fifo_FPGA_to_HPS_out_csr_read                 => mm_interconnect_1_fifo_fpga_to_hps_out_csr_read,           --                                        .read
			fifo_FPGA_to_HPS_out_csr_readdata             => mm_interconnect_1_fifo_fpga_to_hps_out_csr_readdata,       --                                        .readdata
			fifo_FPGA_to_HPS_out_csr_writedata            => mm_interconnect_1_fifo_fpga_to_hps_out_csr_writedata,      --                                        .writedata
			fifo_HPS_to_FPGA_in_write                     => mm_interconnect_1_fifo_hps_to_fpga_in_write,               --                     fifo_HPS_to_FPGA_in.write
			fifo_HPS_to_FPGA_in_writedata                 => mm_interconnect_1_fifo_hps_to_fpga_in_writedata,           --                                        .writedata
			fifo_HPS_to_FPGA_in_waitrequest               => mm_interconnect_1_fifo_hps_to_fpga_in_waitrequest,         --                                        .waitrequest
			fifo_HPS_to_FPGA_in_csr_address               => mm_interconnect_1_fifo_hps_to_fpga_in_csr_address,         --                 fifo_HPS_to_FPGA_in_csr.address
			fifo_HPS_to_FPGA_in_csr_write                 => mm_interconnect_1_fifo_hps_to_fpga_in_csr_write,           --                                        .write
			fifo_HPS_to_FPGA_in_csr_read                  => mm_interconnect_1_fifo_hps_to_fpga_in_csr_read,            --                                        .read
			fifo_HPS_to_FPGA_in_csr_readdata              => mm_interconnect_1_fifo_hps_to_fpga_in_csr_readdata,        --                                        .readdata
			fifo_HPS_to_FPGA_in_csr_writedata             => mm_interconnect_1_fifo_hps_to_fpga_in_csr_writedata,       --                                        .writedata
			led_pio_s1_address                            => mm_interconnect_1_led_pio_s1_address,                      --                              led_pio_s1.address
			led_pio_s1_write                              => mm_interconnect_1_led_pio_s1_write,                        --                                        .write
			led_pio_s1_readdata                           => mm_interconnect_1_led_pio_s1_readdata,                     --                                        .readdata
			led_pio_s1_writedata                          => mm_interconnect_1_led_pio_s1_writedata,                    --                                        .writedata
			led_pio_s1_chipselect                         => mm_interconnect_1_led_pio_s1_chipselect,                   --                                        .chipselect
			RegAddr_pio_s1_address                        => mm_interconnect_1_regaddr_pio_s1_address,                  --                          RegAddr_pio_s1.address
			RegAddr_pio_s1_write                          => mm_interconnect_1_regaddr_pio_s1_write,                    --                                        .write
			RegAddr_pio_s1_readdata                       => mm_interconnect_1_regaddr_pio_s1_readdata,                 --                                        .readdata
			RegAddr_pio_s1_writedata                      => mm_interconnect_1_regaddr_pio_s1_writedata,                --                                        .writedata
			RegAddr_pio_s1_chipselect                     => mm_interconnect_1_regaddr_pio_s1_chipselect,               --                                        .chipselect
			RegContent_pio_s1_address                     => mm_interconnect_1_regcontent_pio_s1_address,               --                       RegContent_pio_s1.address
			RegContent_pio_s1_readdata                    => mm_interconnect_1_regcontent_pio_s1_readdata,              --                                        .readdata
			sysid_qsys_control_slave_address              => mm_interconnect_1_sysid_qsys_control_slave_address,        --                sysid_qsys_control_slave.address
			sysid_qsys_control_slave_readdata             => mm_interconnect_1_sysid_qsys_control_slave_readdata        --                                        .readdata
		);

	irq_mapper : component soc_system_irq_mapper
		port map (
			clk           => open,                     --       clk.clk
			reset         => open,                     -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq, -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq, -- receiver1.irq
			sender_irq    => hps_0_f2h_irq0_irq        --    sender.irq
		);

	irq_mapper_001 : component soc_system_irq_mapper_001
		port map (
			clk        => open,               --       clk.clk
			reset      => open,               -- clk_reset.reset
			sender_irq => hps_0_f2h_irq1_irq  --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_0_h2f_reset_reset_n_ports_inv,  -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	hps_0_h2f_reset_reset_n_ports_inv <= not hps_0_h2f_reset_reset;

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_1_button_pio_s1_write_ports_inv <= not mm_interconnect_1_button_pio_s1_write;

	mm_interconnect_1_dipsw_pio_s1_write_ports_inv <= not mm_interconnect_1_dipsw_pio_s1_write;

	mm_interconnect_1_led_pio_s1_write_ports_inv <= not mm_interconnect_1_led_pio_s1_write;

	mm_interconnect_1_regaddr_pio_s1_write_ports_inv <= not mm_interconnect_1_regaddr_pio_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	hps_0_h2f_reset_reset_n <= hps_0_h2f_reset_reset;

end architecture rtl; -- of soc_system
